//`include "testbench_top.sv"
//`include "basic_test.sv" 