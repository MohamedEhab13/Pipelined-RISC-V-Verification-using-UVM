`include "risc_top.sv"
`include "risc_v.sv"
`include "data_mem.sv"
`include "controller.sv"
`include "hazard_unit.sv"
`include "data_path.sv"
`include "reg_file.sv"
`include "alu.sv"
`include "extend.sv"
`include "main_decoder.sv"
`include "alu_decoder.sv"
`include "c_dec_ex.sv"
`include "c_ex_mem.sv"
`include "c_mem_wr.sv"
`include "d_dec_ex.sv"
`include "d_ex_mem.sv"
`include "d_mem_wr.sv"
`include "d_fetch_dec.sv"
`include "adder.sv"
`include "flopenr.sv"
`include "flopr.sv"
`include "mux2.sv"
`include "mux3.sv"
`include "mux4.sv"



